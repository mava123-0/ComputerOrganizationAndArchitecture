module andgate(a,b,y);
input a,b;
output y;
and(y,a,b);
endmodule