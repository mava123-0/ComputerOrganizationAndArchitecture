module demux14tb_24_05;
reg d,s0,s1;
wire o1,o2,o3,o4,nots0,nots1;
